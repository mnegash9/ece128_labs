module subtracter(input clk, input [3:0] a, b, output [7:0] difference);

    assign difference = a - b;


endmodule